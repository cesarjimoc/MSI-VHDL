library ieee; -- Importa la librería estándar IEEE
use ieee.std_logic_1164.all; -- Importa el paquete std_logic_1164

-- Importa la librería estándar IEEE y el paquete para señales std_logic.

entity MSS_sl is -- Define la entidad para la máquina de estados secuencial con carga
	port(
		resetn,clk,start,enter: in std_logic; -- Entradas: resetn, clk, start, enter
		est: out std_logic_vector(3 downto 0); -- Salida de estado
		e0,e1,e2,fin,resetnReg: out std_logic); -- Salidas de indicadores y control
end MSS_sl; -- Fin de la declaración de la entidad

-- Entidad MSS_sl: máquina de estados secuencial con carga. Entradas: resetn, clk, start, enter. Salidas: est, e0, e1, e2, fin, resetnReg.

architecture solve of MSS_sl is -- Arquitectura principal
	-- Signals,Constants,Variables,Components -- Aquí se pueden declarar señales, constantes, variables, componentes
	type estado is (s0,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12); -- Tipo de datos para los estados
	signal y: estado; -- Señal para almacenar el estado actual
	begin
	--Process #1: Next state decoder and state memory -- Proceso para decodificar el siguiente estado y almacenar el estado actual
	process(resetn,clk) -- Proceso sensible a resetn y clk
	--Sequential programming -- Programación secuencial
		begin
			if resetn = '0' then y<= s0; -- Si resetn está activo, estado inicial s0
			elsif (clk'event and clk = '1') then -- Flanco de subida del reloj
				case y is -- Decodificación de estados
					when s0 => 
							if start='0' then y <= s0; -- Permanece en s0
							else y <= s1; end if; -- Va a s1
					when s1 => 
							if start='1' then y <= s1; -- Permanece en s1
							else y <= s2; end if; -- Va a s2
					when s2 => 
							if enter='0' then y <= s2; -- Permanece en s2
							else y <= s3; end if; -- Va a s3
					when s3 => 
							if enter='1' then y <= s3; -- Permanece en s3
							else y <= s4; end if; -- Va a s4
					when s4 => y <= s5; -- Va a s5, Output Decoder, e0=1
					when s5 => 
							if enter='0' then y <= s5; -- Permanece en s5
							else y <= s6; end if; -- Va a s6
					when s6 => 
							if enter='1' then y <= s6; -- Permanece en s6
							else y <= s7; end if; -- Va a s7
					when s7 => y <= s8; -- Va a s8, Output Decoder, e1=1
					when s8 => 
							if enter='0' then y <= s8; -- Permanece en s8
							else y <= s9; end if; -- Va a s9
					when s9 => 
							if enter='1' then y <= s9; -- Permanece en s9
							library ieee; -- Importa la librería estándar IEEE
							use ieee.std_logic_1164.all; -- Importa el paquete std_logic_1164
							entity MSS_sl is -- Define la entidad para la máquina de estados secuencial con carga
							if start='1' then y <= s12; -- Permanece en s12
									resetn,clk,start,enter: in std_logic; -- Entradas: resetn, clk, start, enter
				end case;
									e0,e1,e2,fin,resetnReg: out std_logic); -- Salidas de indicadores y control
							end MSS_sl; -- Fin de la declaración de la entidad
							architecture solve of MSS_sl is -- Arquitectura principal
			case y is -- Decodificación de salidas
								type estado is (s0,s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12); -- Tipo de datos para los estados
				when s1 => est<="0001"; -- Estado s1
							    -- Aqu ed se pueden declarar se f1ales, constantes, variables, componentes
							    signal y: estado; -- Se f1al para almacenar el estado actual
							    begin
							    -- Proceso para decodificar el siguiente estado y almacenar el estado actual
							    process(resetn,clk) -- Proceso sensible a resetn y clk
							        begin
							            if resetn = '0' then y<= s0; -- Si resetn est e1 activo, estado inicial s0
							            elsif (clk'event and clk = '1') then -- Flanco de subida del reloj
							                case y is -- Decodificaci f3n de estados
							                    when s0 => 
							                        if start='0' then y <= s0; -- Permanece en s0
							                        else y <= s1; end if; -- Va a s1
							                    when s1 => 
							                        if start='1' then y <= s1; -- Permanece en s1
							                        else y <= s2; end if; -- Va a s2
							                    when s2 => 
							                        if enter='0' then y <= s2; -- Permanece en s2
							                        else y <= s3; end if; -- Va a s3
							                    when s3 => 
							                        if enter='1' then y <= s3; -- Permanece en s3
							                        else y <= s4; end if; -- Va a s4
							                    when s4 => y <= s5; -- Va a s5, Output Decoder, e0=1
							                    when s5 => 
							                        if enter='0' then y <= s5; -- Permanece en s5
							                        else y <= s6; end if; -- Va a s6
							                    when s6 => 
							                        if enter='1' then y <= s6; -- Permanece en s6
							                        else y <= s7; end if; -- Va a s7
							                    when s7 => y <= s8; -- Va a s8, Output Decoder, e1=1
							                    when s8 => 
							                        if enter='0' then y <= s8; -- Permanece en s8
							                        else y <= s9; end if; -- Va a s9
							                    when s9 => 
							                        if enter='1' then y <= s9; -- Permanece en s9
							                        else y <= s10; end if; -- Va a s10
							                    when s10 => y <= s11; -- Va a s11, Output Decoder, e2=1
							                    when s11 => 
							                        if start='0' then y <= s11; -- Permanece en s11
							                        else y <= s12; end if; -- Va a s12
							                    when s12 => 
							                        if start='1' then y <= s12; -- Permanece en s12
							                        else y <= s0; end if; -- Va a s0
							                end case;
							            end if;
							    end process; -- Fin del proceso de estados
							    -- Proceso para decodificar las salidas
							    process(y) -- Proceso sensible al estado actual
							        begin
							            case y is -- Decodificaci f3n de salidas
							                when s0 => est<="0000"; -- Estado s0
							                when s1 => est<="0001"; -- Estado s1
							                when s2 => est<="0010"; -- Estado s2
							                when s3 => est<="0011"; -- Estado s3
							                when s4 => est<="0100";-- Estado s4, Output Decoder, e0=1
							                when s5 => est<="0101"; -- Estado s5
							                when s6 => est<="0110"; -- Estado s6
							                when s7 => est<="0111";-- Estado s7, Output Decoder, e1=1
							                when s8 => est<="1000"; -- Estado s8
							                when s9 => est<="1001"; -- Estado s9
							                when s10 => est<="1010";-- Estado s10, Output Decoder, e2=1
							                when s11 => est<="1011"; -- Estado s11
							                when s12 => est<="1100"; -- Estado s12
							            end case;
							    end process; -- Fin del proceso de salidas
							    -- Decodificador de salidas
							    e0<= '1' when y=s4 else '0'; -- Indicador de estado e0
							    e1<= '1' when y=s7 else '0'; -- Indicador de estado e1
							    e2<= '1' when y=s10 else '0'; -- Indicador de estado e2
							    fin<= '1' when (y=S11) or (y=s12) else '0'; -- Indicador de finalización
							    resetnReg <= '0' when y=s0 else '1'; -- Señal de reset para el registro
							    -- Aquí podrían ir más procesos
							end solve; -- Fin de la arquitectura

							-- type estado: define los estados posibles.
							-- signal y: almacena el estado actual.
							-- process(resetn,clk): decodifica el siguiente estado y almacena el estado actual.
							-- process(y): decodifica las salidas según el estado actual.
							-- e0, e1, e2: indicadores de estado.
							-- fin: indica finalización.
							-- resetnReg: señal de reset para el registro.
